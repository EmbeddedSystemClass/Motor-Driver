*SRC=BZT52C15;DI_BZT52C15;Diodes;Zener 10V-50V; 15.0V  0.500W   Diodes Inc.
-
*SYM=HZEN
.SUBCKT DI_BZT52C15  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 12.7
.MODEL DF D ( IS=13.7p RS=31.9 N=1.10
+ CJO=32.7p VJ=1.00 M=0.330 TT=50.1n )
.MODEL DR D ( IS=2.75f RS=14.5 N=3.00).ENDS
