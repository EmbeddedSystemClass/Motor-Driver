* TLV6741 - Rev. B
* Created by Ramon Jimenez, Collin Wells; October 05, 2017
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2017 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt TLV6741 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID 0
I_B         38 MID 10P
V_GRp       58 MID 110
V_GRn       59 MID -110
V_ISCp      52 MID 57
V_ISCn      53 MID -57
V_ORn       47 VCLP -1
V11         57 46 0
V_ORp       45 VCLP 1
V12         56 44 0
V4          26 OUT 0
VCM_MIN     80 VEE_B 0
VCM_MAX     81 VCC_B -1.2
I_Q         VCC VEE 850U
V_OS        39 36 129.856U
C_DIFF      ESDp ESDn 6P  
GVCCS4      22 MID 21 MID  -1U
R73         MID 22 R_NOISELESS 1MEG 
C25         22 MID  3.18000000000000E-0016  
XU4         23 MID MID CLAMP VCCS_LIM_2_0
XU3         24 25 MID 23 VCCS_LIM_1_0
G_Aol_Zo    27 MID CL_CLAMP 26  -89
XVCVS_LIM_1 28 MID 29 MID VCVS_LIM_1_0
R70         28 30 R_NOISELESS 10K 
R61         28 MID R_NOISELESS 30.09 
C23         30 28 53.05F  
GVCCS3      30 MID 31 MID  -24.6
R57         30 MID R_NOISELESS 1 
Rdc         27 MID R_NOISELESS 1 
Rx          26 29 R_NOISELESS 330K 
Rdummy      MID 26 R_NOISELESS 33K 
R55         31 27 R_NOISELESS 10K 
R54         31 MID R_NOISELESS 66.67K 
C21         27 31 79.58N  
R65         MID 32 R_NOISELESS 680.9 
C22         32 33 99.47P  
R66         33 32 R_NOISELESS 10K 
GVCCS2      33 MID 34 MID  -15.69
R69         MID 33 R_NOISELESS 1 
R64         MID 34 R_NOISELESS 1.997K 
C20         34 35 31.76P  
R63         35 34 R_NOISELESS 100MEG 
G_adjust    35 MID ESDp MID  -1.5M
Rsrc        MID 35 R_NOISELESS 1 
C15         21 MID 8F  
R56         MID 21 R_NOISELESS 1MEG 
GVCCS1      21 MID VSENSE MID  -1U
R44         MID 23 R_NOISELESS 1MEG 
R68         MID CLAMP R_NOISELESS 1MEG 
C36         CLAMP MID 2.3N  
XIn11       ESDn MID FEMT_0
Xi_n        MID 36 FEMT_0
Xe_n        37 36 VNSE_0
R51         ESDp 37 R_NOISELESS 1M 
XVOS_VCM    38 39 VCC VEE VOS_SRC_0
S5          VEE ESDp VEE ESDp  S_VSWITCH_1
S4          VEE ESDn VEE ESDn  S_VSWITCH_2
S2          ESDn VCC ESDn VCC  S_VSWITCH_3
S3          ESDp VCC ESDp VCC  S_VSWITCH_4
C28         40 MID 1P  
R72         41 40 R_NOISELESS 100 
C27         42 MID 1P  
R71         43 42 R_NOISELESS 100 
R75         MID 44 R_NOISELESS 1 
G14         44 MID 45 MID  -1
R74         46 MID R_NOISELESS 1 
G13         46 MID 47 MID  -1
R46         MID 48 R_NOISELESS 2.083K 
C14         48 49 63.66P  
R48         49 48 R_NOISELESS 100MEG 
G6          49 MID VEE_B MID  -67.6M
Rsrc1       MID 49 R_NOISELESS 1 
R49         MID 50 R_NOISELESS 2.083K 
C16         50 51 63.66P  
R50         51 50 R_NOISELESS 100MEG 
G9          51 MID VCC_B MID  -67.6M
Rsrc2       MID 51 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
XCL_AMP     52 53 VIMON MID 54 55 CLAMP_AMP_LO_0
S8          CLAMP 56 CLAMP 56  S_VSWITCH_5
S9          57 CLAMP 57 CLAMP  S_VSWITCH_6
XGR_AMP     58 59 60 MID 61 62 CLAMP_AMP_HI_0
R39         58 MID R_NOISELESS 1T 
R37         59 MID R_NOISELESS 1T 
R42         VSENSE 60 R_NOISELESS 1M 
C19         60 MID 1F  
R38         61 MID R_NOISELESS 1 
R36         MID 62 R_NOISELESS 1 
R40         61 63 R_NOISELESS 1M 
R41         62 64 R_NOISELESS 1M 
C17         63 MID 1F  
C18         MID 64 1F  
XGR_SRC     63 64 CLAMP MID VCCS_LIM_GR_0
R21         54 MID R_NOISELESS 1 
R20         MID 55 R_NOISELESS 1 
R29         54 65 R_NOISELESS 1M 
R30         55 66 R_NOISELESS 1M 
C9          65 MID 1F  
C8          MID 66 1F  
XCL_SRC     65 66 CL_CLAMP MID VCCS_LIM_4_0
R22         52 MID R_NOISELESS 1T 
R19         MID 53 R_NOISELESS 1T 
XCLAWp      VIMON MID 67 VCC_B VCCS_LIM_CLAWP_0
XCLAWn      MID VIMON VEE_B 68 VCCS_LIM_CLAWN_0
R12         67 VCC_B R_NOISELESS 1K 
R16         67 69 R_NOISELESS 1M 
R13         VEE_B 68 R_NOISELESS 1K 
R17         70 68 R_NOISELESS 1M 
C6          70 MID 1F  
C5          MID 69 1F  
G2          VCC_CLP MID 69 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 70 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 71 72 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         71 MID R_NOISELESS 1 
R24         MID 72 R_NOISELESS 1 
R27         71 73 R_NOISELESS 1M 
R28         72 74 R_NOISELESS 1M 
C11         73 MID 1F  
C10         MID 74 1F  
XCLAW_SRC   73 74 CLAW_CLAMP MID VCCS_LIM_3_0
H2          43 MID V11 -1
H3          41 MID V12 1
C12         SW_OL MID 1N  
R32         75 SW_OL R_NOISELESS 100 
R31         75 MID R_NOISELESS 1 
XOL_SENSE   MID 75 42 40 OL_SENSE_0
S1          27 31 SW_OL MID  S_VSWITCH_7
H1          76 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_8
S6          OUT VCC OUT VCC  S_VSWITCH_9
R11         MID 77 R_NOISELESS 1T 
R18         77 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 1P  
E5          77 MID OUT MID  1
C13         VIMON MID 1P  
R33         76 VIMON R_NOISELESS 100 
R10         MID 76 R_NOISELESS 1T 
R47         78 VCLP R_NOISELESS 100 
C24         VCLP MID 100P  
E4          78 MID CL_CLAMP MID  1
R62         MID CL_CLAMP R_NOISELESS 1K 
G4          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 22 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          24 MID 1F  
R9          24 79 R_NOISELESS 1M 
R7          MID 80 R_NOISELESS 1T 
R6          81 MID R_NOISELESS 1T 
R8          MID 79 R_NOISELESS 1 
XVCM_CLAMP  82 MID 79 MID 81 80 VCCS_EXT_LIM_0
E1          MID 0 83 0  1
R77         VEE_B 0 R_NOISELESS 1 
R5          84 VEE_B R_NOISELESS 1M 
C3          84 0 1F  
R60         83 84 R_NOISELESS 1MEG 
C1          83 0 1  
R3          83 0 R_NOISELESS 1T 
R59         85 83 R_NOISELESS 1MEG 
C2          85 0 1F  
R4          VCC_B 85 R_NOISELESS 1M 
R76         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R67         86 82 R_NOISELESS 1K 
G1          82 86 50 48  -1M
R2          25 ESDn R_NOISELESS 1M 
R1          86 87 R_NOISELESS 1M 
R58         38 87 R_NOISELESS 1K 
G5          87 38 32 MID  -1M
C_CMn       ESDn MID 6P  
C_CMp       MID ESDp 6P  
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_8 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_9 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

.ENDS TLV6741
*
.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1.65E-3
.PARAM IPOS = 0.247
.PARAM INEG = -0.247
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCVS_LIM_1_0  VC+ VC- VOUT+ VOUT-
.PARAM GAIN = 3.333E2
.PARAM VPOS = 1E6
.PARAM VNEG = -1E6
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=2
.PARAM NVRF=2
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=100
.PARAM NLF=8
.PARAM NVR=4.5
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VOS_SRC_0  V+ V- REF+ REF-
E1 V+ 1 TABLE {(V(REF+, V-))} =
+(0, 1.6E-3)
+(1, 1.6E-3)
+(1.3, 0)
+(5.5, 0)
E2 1 V- TABLE {(V(V-, REF-))}=
+(-0.7, -2E-4)
+(-0.5, -2E-4)
+(-0.4, 0)
+(5.5, 0)
.ENDS VOS_SRC_0 
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.035
.PARAM INEG = -0.035
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.440
.PARAM INEG = -0.440
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAWP_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 5E-5)
+(10, 1.38E-4 )
+(20, 2.93E-4)
+(30, 4.78E-4)
+(40, 7.21E-4)
+(45, 8.95E-4)
+(47, 9.92E-4)
+(50, 1.24E-3)
+(52, 1.59E-3)
+(54, 2.23E-3)
.ENDS VCCS_LIM_CLAWP_0 
*


.SUBCKT VCCS_LIM_CLAWN_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 5E-5 )
+(10, 1.29E-4)
+(20, 2.77E-4)
+(30, 4.52E-4)
+(40, 6.77E-4)
+(45, 8.31E-4)
+(47, 9.09E-4)
+(50, 1.08E-3)
+(52, 1.3E-3)
+(54, 2.25E-3)
.ENDS VCCS_LIM_CLAWN_0 
*


.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 220E-3
.PARAM INEG = -220E-3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIM_3_0 
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


